PK   qGVFV�tT  �J    cirkitFile.json�]ے�6����&V��K��g��3v�'��
^݊UK���m��?h~f�iJ��H�<��rtu;\�B"���d��6��\/�Ͷ\�Znw��zv��|�1����߲��a�^�7�_�������s�����ͧ�ͺ\�R�i�D�aT*�Y�i�,��GYT�����uu�R�"̓X�<P���DK�L	�
�H���/�;F.R��L'A�U��� �b��yTeEQ�O(C�Cs���1r�LJ��,e�d���C�Q�a"�,�*���vӭ�Є�C��y�$HD��Ȣ �X�
)�L�J��,r��IX%3�Y��LW"�0ETe���*h#ǎ�9y��,Hd��
�q�L�B��&>s��ʲ�̩��8M��l3c1��L�*R�X��8PI^��a���R��D�Z�sZwA�.i���{�Aݝ;,W"DEf��`igY�i*T��,s�! ��wm�R��v�h�H�����$U*ˋ*(un�����a�y���(,�R���MƉ���'�3N�h<$�'��'��Жs�xl�Һ��uwc��2�T��*:���
%93�")���L�w�Zhd7h��n�B�ݐ���u'�SK�l����Aۣ0��D��(L�?}�eaD2��ks�����͆��H���
�YR�]�9rq����̌'2�j�ܞ�:�i�CQ&����X����̌[V�ғ��ޘĢ�%�y�\}��2�G���fV��82ƒXU����ٷ*E��N�Rc[D���"�m��(Γ�p�]nYw_Ȧq���ؽĠJ�t���]�C���'jDAԈ�u��Σ�%�\0���X� *bA��k�����+'ҲI�n���&�63q�I��!���D�K7�!�u�'�>Aۅ�Z�CC��InW�p��!����$�+h�M�А��zh��4�'Yi�Jv=4� ��S<4h��<�݊Q���B	�?��:���i[9����kP�uK��(��[j�	z�4�k�@%D�dvKp�;�&�5x�����'�Ææ�`=:�\d�Ԯ�mGJ��[j0���Ԡ� 5	ׂ�C�K���L�Z"��	b�f[Rf��ݫ��	ft����"�s��#�N�F�����I��"��j�%&Dξ5'��Cr�.<�	\��R�,#�"-Ʋ�U����'�Y���k�K��~"m�O��\83�	�Kb�Ĺ��A�?�h"�.�酋��e�h�]�~A��<��i4�_K�Ym�j
�P������/�`��<����y�M2�Mp��e�h��.�F��fߦ"*uA�2�_4���A���m���.�^?���p�6�N������50�#�o��yX�����Cyz��~P,��X�!S�%�!�?(~T�H��X8������ғ)��ҏ.�~P,��X�������?�
M�����)9����5��4S�_4��c�&�����o��y%���)"��?��ѿ��~YЌ�~ԡ�����+�F��eA���; �n�˂F������h4��<C��Z
�U��1h�_4��/W�R`��F�a��>ݗ԰Ӻ|�o�1�D�"�p�^�(/\�.�.�.�.�8�D�2�]8�D�2�]8�D�2�]8�D�2�]8�D����x�����/��_�����s?�~@�Q���\1���\���\����\����\�`wX�a'l��wX�a'l� xX�a'l��ؓ~P,<�`?(~P,��X�A���b�����K?(�~P,=�~P,��X�A��b9�b8�D�2�8�D�2(v�s�;ѹ�v�s�;ѹ����\e��Nt.���a':�AY��ˠ,p؉�eX��a':�AY��˰~A�Nt.�|����?��X���>/��n�2:�X,׋Ͷ(���w��g?l>��`�.W�"�A����QC:��:QhF�D�rc���U�]�7�w�s_% H���_\����7^.=Ί��r�9(C�K%���:o����"k�b��h�8COSF�CSj;��ʟ��0ń�׃)�olS^�&�M3����R^.�佈\��{i%�|���"HYgG�LЭDYgJe�:S�/;G�<��cd�OqM02\ʊRv��z5��Ա	v\`ɻ&�����sB���aE�����Tp0�U�����~����{�!����Rp)�W�Д�v�k�y��~K_m�)_3�W�|��CSj���b��\uͿ�64��˚z����Շ�Xɶ����,�芛�32⷟o?�~�����`��<�TG��MB��D�H��v��m`}��Wk�D��Jp����9�ϧ[4�>�vEC��I�F�{%�J`���7>�>�*�a��$@���I��'� ��O�D4�+�5"��V�b�\#��+�5"t��t��tP}J}\#t�+�5"��	���ېϟ�hX�m�F�'SDh��Ɩ��NS�"�0�=_�,� <ϼ�f��Z����\##�>�Č�<Fh~�O@�X�@��p�«<��*��x�p���\%}�3.rCG��9���w����8��>Ө8ՆE�7���U���/-��y�kib�}
�Pĝ�x|o��UR��sp���\#%�xu%�����URӌ�t[<.ק�ҧϛ�r���㲠֛f�?��X���L�+P7�QC���qr�5�=>�-� ��Z�P��6;MrK��9�5\���."ԙ{��Ք���_�+b���e�15ק���V�ΆKTcj�U��1�h5	�T�r*~9����(*��u!T��� .?M�߃C��4�
�2Ӎ}IIq�$\i�ҿ�puiJ*9�T@�)F�~4�A�b�kF�Paا�
јu������f4I�'���Sѡ;I�4*l��
[A՟��O���TRq*�'<���O%��
L�L��sVG\���p��7��. �IW�nps�-��Иtpm�7��.�Z-������J׏npsp!�;�&�+Jc����1�5�1��b�P�Әtp��;�&��Pc������L�`G�f�7W�	�U�I�nps�[p�jL:��5&\��.l�Z�/��3�ea�]�����(������d!b���D-�햳*�*[�e���p���&��ܒrK�-1��ܒsK_���2�3�|�R���5o�C���������=��Q��H�C��������=��!m��b>?�逘g��b�\� �����r�^t@ċ�u�96.: ��r �z��w�� ���F�<�ͺ�[m�0��M}wߙ! ^,(ᲗGNi	Քk嬡���Ŷ�\�(�ZT�܁rJn��)�-��5��2��WJ�0h/R,aZZnk
�c
)o�Pj��P��"ʕ��� F(
�����@��xn(9\��+��!��s��A�ôWb).���D�3�(n7��� ��A��8%���>��/�Z�Y��fz�>����cGk5uo7�c�h7�c�l7�c�j7�c�n7�Ǧ����vS|l���$]�ٶL�l�nm��j�X-w{��P��P.��_������UY��n7�g���ҽ�f�Q�������e�����?��aw��r��y�u��~���ٯ���~2*�|z\/� 3������5<g�U�ڕ�qWn^�٪<�n[���r[����of�S�~��|���u;݃��=K�f�n��o�_���y�TF���n�_n�|�d��<G�\��.IB��D�̱�{�c��'
��t�����T�R�*�B�#�r�ۧ�����g��}zm��`~�/���<.��6wz��an>��N�z�c#p(œı�U7=�{��i�X,7?��݁)��ẁ�!0B�bw�oT@�4\ �C]��KaQq�31-��C"��?j'�+T�@�T*��Sg�&ќ3�kਨ	Ӥސ3�٣�%r找��r�C'�9l.���ܰ��!��8��7��F�n�&V��ɚ	� �2ji��i�hQ��}��X-P��9��oYF�'�.�;3� K*y�y�U��y�+��Ny��<�l�
�"`���K1��͙(�\-���:��v��"�}���n��㑩�-a|G5�	�c�'ԝ�39�e5��3��1uq�jk�X����̺�Y�!/� �xl��6�WQ�TU��;�� �a�6�O��G���yy��Ly:]OML4�wlJ��)����%{C��;����RS�����Aؖ�Aؖ����Y���O�M'����ڍ�i\ޙ�I��A���N�Pq�]F�HG:fG-ᢋ�;��X�㤛k���D���D��D<c�Ihǌ�
��|^;��BI7�z"�^x����-��L%�G�gO*���0fu��Q�߿J����~�{/���_l�
�'f����v)�$ܺ#��Y�ۦDF�b�y�,�3ճH�/v?��S�D�+v�?�O������#��u�u诖��㧬�~�C��w����פ=��BH57�|h���Ö� ;W���#m�\��2`�����,���ѕq�[�ʲ��:�k��u�ږ7�~]���1�Pذ��Dz�$z��̯���u�d`B�~0�^␋�Oo����ilŻs����#M�)�a��4n������-o����[��Ȁ�2�!���&e��z:|z�WL΄dB����)<�f�A�k��b^Ny����8�������4d�i�JE�AA�cA7(U��\�Ö�j[^��4�^c��N�v]LC�*)�*��Y��R:7�¢�����6�9Ы�cbJ=�.�?�_���p�S����n�ι'���S��������[�p�ĉ�O;�4 ���v���q��s��QTGK���"��{���:�+� l�{'a
��"�T�k㥛���n�6�:�:��M��Y7]u�tmvӵ�M��g7]��t��k#�M�f7|]v�ti����o�lе��E2fC��bٖ!�������Lo��̄���"�~G�~X���m6G�����)�]~��\����re4V�u��Z����}H�e���%���~���������A��{��V������ٷUe�������L�v��r�}Q7����Y�.zY���ּ���|�f���G�6����t��f�����g����m�Ou���������鍀�ѷxz/���R̻�Bv~&����Fɬa�Iw���E������=����o����G���'���y[@jЉ�JwS(a5#n���J��QN�Fu��&Yؽ�*bg�Gɸpеp	���X����r�l�ƥ�8Oo���٠��Jw[(A�Kn%\�C��:�	"�J-�-uv�ƗK��IB��)4��I4�BJ82G� s�tc�y�V��9������"�h��1C�U��~��~�tc~x��T8�xu�C/���>׿��B�-����M���١ ŋ�nz�`�� �aU�pč@��F�L9N��=�3K�Ev3��1�SH#�n$XyD$�@7�ҍ��J9�ԥ��M���~Ĕ\�L��޵��j��7	_��T�,�{���>��|�}���>!v�iсGȨ�^ԈP�/5~�,G��K�8C�tBv�%��Z��j��3EG����2E_�������MB�9®�FL����80�R= k�X�[)Ʋ�U>�x�!�ߋ��T�e1	��hҹ�$2X=,=VXܟKԷ=(��D_h^��t����~�|�9|��!����Ж޹T�%Վ0H�B�)�����w��"�jܡ�o�ۿ>-�أkDF��͉�2�<�R��r_.8�o:��M����7oj:�p
|b��q|�����lz&�N�Nw{D�F6J�'��+���n��M�ϱ��w�`ζQk�l���8�p��.}�B-��t-�\�Q���Q�b�K0����9��fH���a�����Fk��)w�hK��t--����[-��&[���:�yXx�+�n��#D��«Ƃ*pAQ:p�+]2���z4Gx�G���|�g]^�d�t����2��i
\�����Q���!�&�!�m�q��	=�b����£t�}Bg��;�M� !�/S�Y�6}�����Gɜ�ͺ n/�x`_�zx�������h�9�?���� ��l=�7���}����!�X��f�q�hҹ�(���3�����˕o��M�_Fg�>�G,<��������8t�t����B���&�#���nz	zu�+�o��� ��)�o�7�\Ϊ�.|*�R>�Uؑ�}3�gg|$��n��bN(��R�t�H��6m��u�"��&���M�&����L�L����z��������.��nvo1��?,��,�����w�O���O;�`�̾�?PK   qGVFV�tT  �J            ��    cirkitFile.jsonPK      =   �    
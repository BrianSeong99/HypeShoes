PK   �qiV��  �n    cirkitFile.json�]�r�F�~s#�?���ك3v�'���@ nƪI-E��u����3mII�>0�<���m	Y�D�WYY�Y�̶ٯ�z��l�ů��a�Y�n���>f��sv��p>�_����mv�qv���9��~_�ͧ�ͺ\�J&Y�e�Q\:[�A^dU �DI�q�L���ݹ�2�i��U��J�.� 7&
D��t.�8Ur�����*SJ�*(�(�H� �c�B�2/�	�r!η�*��ef_ڶey�A�&��H�R��f��(싢0
�̭̙<Z�Hd��d����yU���Z�N�e�I\:�DWaY��mU�e�A�3�
�4�]-�<��e���6�FIxF	j��K�pB�Zz���R%2[���K��U�F� ��0��5�����Y��J)'U�@�TiE�GSF�t�Q�ެ=oN���"��ts��-�El�0%�\�J��H�Ajc�&4�(�T�	){���4��<������V�"
dWE��2�
��"I�x�a$��ʃT�V	��	���Uf�_)��x�R�$�S��U����,��SWVخ��0	�Un*���Ii��;-���\Қ+ZsMk��(�eAP�5J�KL�h�����Yh�ܤA�Wvjk����M'�X�U^U�)�}s;Yj�Ei�En�yfA��Q�e��qR�v�z�-l����4�:aY���,�2T2�=9�V�(��]�����-��[�� �oA��""�'�5�ۧ��Д�/-،�5��j����g#륩�\���+�����++!����̧�!�������5��j�G;ԜvAE;��kO|�����סl��D�	�eyH�V����S�D�K��'�^Q/}z����^M�0�8a$q�H���>ԓ`�m@D�"�^Qm"�Q�+"t��]�%G��F�}���#�9��y�ok�7��`f�o]��7�l	0j5�8c{��owz�7���`��x}�RFм����_PL��_�3�7�`Xa�M�������0��a�S��f#h|����@�&����d��|�A!_���\B�I�Ԕx��i0<G�x�	R�J��S�� �?�kB`�3P BR�
�(R �ް�"�H)�L�����y�Q����,���n�%fAξ��m����e������E:.e��$Y���yV�����,�ލ�cdJ�x�E�"��%�saXQz7u\������ݻh���E�p�,\z���3u�4��A��oN�I?�Z
N��VSp2����������A��x��`X$<l�>6h.�^��=\z���̾�d\�����h��^���8\x�+��˃�~��p����p��k`8��ۤ��s��8ՆCy2�`KK�g��)5��X�X�b����p���̓b�dJ�X��bŃbŃbՋb4��3���t+t4�ۿ���t˂��t�W�t�nY�ԑn����/`JG�]��gt˂�Zt��h�C�@��eA�
�Q��t˂���G�w˂�һg �Swk)4��=�p�y�U{���cиa�,h�[4�֣��0�����vٮ������n���Nt.���b�Y�.���K��%�����\z����\z����\z����\z����\x�+��˃^�_��_�`��`�a��a�bыb8�D�ҋa8�D�ҋ`8�D�ҋ_8�D�ҋ^8�D��~�������_�a'6<���x؉���4��A�d��<(�<(�<(�<(�<(�<(�<(�<(V<(V<(VL�����U/���K/j��K�,p؉ΥW8�D���/h؉ΥW8�D��+v�s�;ѹ�����\ze��Nt.���a':�~�����\ze��Nt.��;ѹ���en������bU�6��|�y�-�wVg��z���vv���,���s����nQD.�������j�䁕�2���+��Kk��7w�v���6~�}�DI�DY���D~]�pI�b��ae�;(��������Ք#��1X�W{*���1z����3��5���_(W���J|�np�n�x5�c���m�W��D�an�<���K����p�|#
��F��5���(A�8Skz\�.{m�J���:1'�m�y�$�q���Ǌ�	|k;�໨�g|��&�ﴻ�5���b5�b�(�8ϛ)���w$����;��/Xb�n.S��\��}4�
�;���|e���6��$ek�V�I.d�A
���~�|�����I*^�
 �Ģ�P�@_�6���+��4{��X�\��I�^�ֻfP*"���*�p1��נ�`K3��h^��#x_A_��Wп5�]��F�K@?��W�˄��@y3-XHy3-BJy3-JIz3��𔟴-?m~-�E�.��*��2Zⷿ��~�����߯'��A"�<�A}v��ƽD�H~\�z�}rX����c��)��L����Ԅ���[o��>��$@}k�L���^�����t�6��u<	�-��[�ѐ���vJ0E�k��7A^Q� S�u
0E���X:�	�t㸝L�.�)�Y��	�&�ҧ!1�v4����MC4�v4E�&�^�2�]�i�R/�]��I��.���E�7���Z$S�?w
0E4���Уy��	����%L��!�W��|�*�lص ����������\ё��'�&���ML�N�$�~� �rѡ�Y�K@Z��)mݛ�)�е4�����ę��|�eb���>����S� n]�.����8H��0�BQ/�-Gʡ��*�fc��la�8��
c��A����d��H�P�S[��<�	0���6�,i'S���7є�7���3-�8jFT#���DV��t06Lq�. ���+I��3�SG$��cw�����8�^�7��wJ�d��0�AQ��D�G�z�x`u?
������Y���Q}iS�%faP��8v�ă���{Gt߀�#J fy��D�2�G�`���bS�lM ��S�sM ��
��z�̲m�Z?׈�yS�ٻ򏫂Z>>l�!�p[�<pA�;JΩj�������-H�-q(Ί��ΐ2�[�(Nƴ��c�Õ�=}נ�������^�w`�2��!��<E�3`��l��<������kГ�O����WP,���8&1��v_ט� �3���S�w�� Oi߁B�j|c^R�����S�w .OiO�� �
�.ň��'1�P�x	x*�#^��.���y���'�=���TRq*��NRt�
[I����VR��<�SJ���TQq��+<���O��
L�L�h{VG\���p�7����Ivop��-�
�tp��7�����Z����v#*\���c�u��<�.�IW��`��Ǥ�k�c@���c�����|IhYyL:��|��G}��(9�g���b���5��<�\���J�I��Ǥ��ԷF��|��fU�x����^H�`v�n�drq���S��n�9��������p��fO�(�#�V8bᨅ#�~�a_a��oc�`9�r�۵����F�ZH�B�ҵ؟�U��r-�^�B�ʵP��r�g�-��q�b�� S�b��� ���R_k����ȂXk��Q�ȲQk�h��8 ʵ� �w�q T�I�w�f]Y؇�M}w˞�3���jN��Q��*J��Plʶ���$���P.<(�\{0��:S���l���������#�q �-�]�<]H���rڅrT�rΈr+�65�9�fxm����<b(������!��!��׼�>$��a�m��h�CbʈxV�Iꗶ�b�?d�`)n��|W��[�eyy����}>�{���閶Q�$ڏ��l?R�G��H��#s|dڏ�㣨�(>>�ۏ���9H���E�-�"�d[W��,�V;7�P�H-�������we��ouϳ�p�y�k�s۬?���q��/��U�w�|�_����Zav����!����=��~���OV�ڟ�+���������?�����V��Ci>�۟W���|�ݶ���ն�{ϝ��ħl�Xe���֕����E��3u���}���xtm�Х�b�oV����ǻ���&Ts�ӛ4�tz��(ۯN��m��Ҫ<Y�Y`��.�N�Bde�Y�ZdERX�V�]�^�@ޕ�lc?k���������<��0�7f�ExSꇹ}�7�$�b�s���|�Ub\�e�_��O��b����>�&n�Mh�.:�� ��;M�6t�ȁ�lrt�㠢#��7�0"EF�Y�BE�SE�!�tH�@G��Qᡌ�ǩ%ӂ
y	���T��P�->O�Qz�����7��F����m�uUA�#t|�Ӛ�G�u �3\��S��|58�¡�叙[[�&r����S�dJ$I����J�@�L��4���H�R�M�@_&2��$��P���52� ��sT^B����r�%�(Gq����>:����(�>�I/atd��n��މ��F��*I�"�-̍�L�j�NF���N@�Bi�*"QfA��$(ef�,��22��Z�9�	LOY[��<�u���b�G ���GW��.<��-��t*=
��n���O�ž��>Ԃ���G5��G��Ta�[=������G����2��p�Md��Q��Z�V���0�B�n:��b�$4>�Xݨ0I�8�Sm��G'��h�p����G�d��vc���Cg�*����G��:���Sl�jx�<'D��H���:j���߆�qj��V��W�?��/.1'��v��V�ckF�¹a���+�M�������E����_���wj�a�zq#��
o���O����?�ÿ8��5�R�����o~���.[��5iO��	��fA�o�GJ7�#����el�:ͳL�.����K�*m�r�4-��a&Q�RT{����Q�7�~e����ABF-����V�MKs���:������2�oȘ�� 1̚�:5�e�u���_6�;�z*�bJ����=6�29�|���_#6�P�� l�:6�6�:l�i�*��<y/��ԽLG�궸o���P+�@k�]
���R��K�gL��ܣKܚ˩���!=�h�׵����ZVQ`�Ƀ�*u`���.
a��Ya����+�A:�W�p?�uz��Q*k?���Q���?U�~z$Z���Ga3z���4�X'Obo�m��mꑨ����5ҩ�E:񶉼mZ!��'���8r�.>�:���a��2�j��Z���C�F������tm�x�Z��еP�ka�C�F������tm�y�ZX�е��k��C�Bm���>��샤����d� :O���	s6������B�I���nny/� �3'^�q���P��Cl�z{s�>+��&�q�����Y����B���yU�>:Qb�~q���r��GGkW q��d���V��O_�.�Ȗ���#?n�����W����c�����ĺ�l��n�Ͼ�*�u�g��3ۭ�ݏ�������G����u��
<����>��)������oV�ݏ�����߿��30?T?�?��}�oo߹���������p4�a�^HX�	�J�	���X>�jg��N�_�ϾX���a�\w�vn�q��6_�"d ɀ��	v_�a��� �� �)<�B�@��	@2���@�]d��@2@:2H�C
�}�0BA�"d 	v��U@2@�+���Ѻ8I5�c�ˀ���Z  �x i&��nu'6.�{y1'D�\D���p��\DH7"�#u~H�'���Ϧ�ad���8�]�v2@�몐��q�8�ϑ�FџN`��]K�����~�%E0��m�Z� ���q����W��Rȫ�����x:a>��G�9/>$��Mf|H����I�ߛ��yݴ�X�9B,a����`i�h\.��T?�۵nz����=��~���z��k�}�,��)x��t�x��
�y�U�	�j&a�'aũ�cЍ[�ިۅs�~�B��oz*M<���A���,�'�k��R�����ƚ��&�Ϗ}�H��|���p� ,�^Sci�b�&��g�ӐJ0��"�*H��U��(�:�$e��wP�zL�����i�	A�E,�? ��B���{��i�h����� QƷ���BB0�2h챂 Xpv�X��� ѐ�,.�����H%��'l��u�=V��Zc?@�ǾA�n<O�06ڄc�ƹ����c/C��!�	�{���U���]{��h���w�WUs��	G1��]H�*Hx�r.t|6G��&��(l�&$XI8>�p�=V�\��T��j�;��,ow-���$A]�$D��)C�4,��;ȼ�������[�{��MB�;�(��q��J����@2@��@{RpLR[E@2��yz��+^|�|�,n%���.U"�%-��� �,>�4�6(!���"+���  ��_]��g&��Y�z��$�t��*B۵�~Qƭ���ƅ��wp�C~�&�7��|E�H8
H�˩nK����"�t���!M��&F�J�Z"ɒX&0V�p&� ���w0���\y]C�� �֐�n�!M<�pY_>@2t�g2.M�Sc���2 ���B��hޤ��5	�2'��[F/!D/q���a@2@�+�DC��Y�<�.j�L7!�܅z�����e�r���f���V�S�֏��w�O���O��>|�}�PK   �qiV��  �n            ��    cirkitFile.jsonPK      =   �    